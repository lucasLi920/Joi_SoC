module wdog_flag_gen #(
  parameter   WDOG_CNT    = 16
) (
  input   logic     pclk,
  input   logic     fclk,
  output  logic     wdog_intrrupt,
  output  logic     wdog_rst_flag
);
  
endmodule